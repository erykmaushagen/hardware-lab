library ieee;
use ieee.std_logic_1164.all;

entity ps_ff_tb is
end ps_ff_tb;

architecture testbench of ps_ff_tb is

--missing

begin
   
--missing
   
end testbench;
