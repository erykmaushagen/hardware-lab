library ieee;
use ieee.std_logic_1164.all;

entity jk_ff_tb is
end jk_ff_tb;

architecture testbench of jk_ff_tb is

component JK_FlipFlop is
    port (
      J,K, clk , reset : in std_logic;
      Q : out std_logic
    );
end component;


--missing

begin

--missing

process begin

--missing
	
	
	
	
	wait;
end process;

end testbench;

