library ieee;
use ieee.std_logic_1164.all;

entity SR_Latch is
    port (
      S,R : in std_logic;
      Q,not_Q : out std_logic
    );
  end SR_Latch;

architecture Behavioral of SR_Latch is

--missing

begin

--missing

end Behavioral;

