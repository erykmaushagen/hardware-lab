library ieee;
use ieee.std_logic_1164.all;

entity ps_ff is
    port (
      d, clk: in std_logic;
      Q, not_Q : out std_logic
    );
  end ps_ff;

architecture behavioral of ps_ff is

--missing

--missing

begin

--missing

end behavioral ;

